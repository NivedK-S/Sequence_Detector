module FSM101Mealy (
    input in,
    input rst,
    input clk,
    output reg out
);
reg [2:0] state;

    
endmodule